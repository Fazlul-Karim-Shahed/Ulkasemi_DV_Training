
`include "apb_interface.sv"
`include "apb_packet.sv"
`include "apb_driver.sv"
`include "apb_monitor.sv"
`include "apb_agent.sv"
`include "apb_scoreboard.sv"
`include "apb_environment.sv"
`include "apb_base_test.sv"
`include "tb_top.sv"
`include "apb_slave_1.vp"