

class apb_packet;

	function new();
		$display("%0t APB Packet constructed", $time);
	endfunction


endclass