
module main;

    int arr[2][3] = {{1,2,3}, {4,5,6}};

    initial begin
        $display("Array: %0p", arr);
    end

endmodule